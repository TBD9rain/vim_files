//  head info

module module_name(

);

//=======================
//  PARAMETER DEFINITIONS
//=======================



//=====================
//  IO PORT DEFINITIONS
//=====================



//======================
//  VARIABLE DEFINITIONS
//======================



//===============
//  DESIGN CODING
//===============



endmodule
