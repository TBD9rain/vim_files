//  head info

module module_name(

);

//======================
//  PARAMETER DEFINITION
//======================



//====================
//  IO PORT DEFINITION
//====================



//=====================
//  VARIABLE DEFINITION
//=====================



//===============
//  DESIGN CODING
//===============



endmodule
