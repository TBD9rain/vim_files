//  head info

module module_name #() ();


//=====================
//  VARIABLE DEFINITION
//=====================



//===============
//  DESIGN CODING
//===============



endmodule
