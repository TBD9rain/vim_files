//  head info

